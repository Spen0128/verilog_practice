module full_adder_4_tb;
    reg [3:0] in_1, in_2;
    wire [3:0] s;
    wire cout;

full_adder_4 main(in_1, in_2, s, cout);

initial 
    begin
        in_1 = 4'b0000; in_2 = 4'b0000;
        #10 in_1 = 4'b0001; in_2 = 4'b0000;
        #10 in_1 = 4'b0001; in_2 = 4'b0001;
        #10 in_1 = 4'b0001; in_2 = 4'b0011;
        #10 in_1 = 4'b0001; in_2 = 4'b0100;
        #10 in_1 = 4'b0001; in_2 = 4'b0101;
        #10 in_1 = 4'b0001; in_2 = 4'b0110;
        #10 in_1 = 4'b0001; in_2 = 4'b0111;
        #10 in_1 = 4'b0001; in_2 = 4'b1001;
        #10 in_1 = 4'b0001; in_2 = 4'b1011;
        #10 in_1 = 4'b0001; in_2 = 4'b1101;
        #10 in_1 = 4'b0001; in_2 = 4'b1110;
        #10 in_1 = 4'b0001; in_2 = 4'b1111;
        #10 in_1 = 4'b0011; in_2 = 4'b0001;
        #10 in_1 = 4'b0011; in_2 = 4'b0010;
        #10 in_1 = 4'b0011; in_2 = 4'b0011;
        #10 in_1 = 4'b0100; in_2 = 4'b0000;
        #10 in_1 = 4'b0100; in_2 = 4'b0110;
        #10 in_1 = 4'b1011; in_2 = 4'b0101;
        #10 $finish;
    end

endmodule
